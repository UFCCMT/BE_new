-----------------------------------------------------------------------------------------------------
-- reg:
-- Description:
-- This is an enable based register. 
-----------------------------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity REG is
  generic (wid   :     positive  := 16;
           init  :     std_logic := '0');
  port(clk       : in  std_logic;
       rst       : in  std_logic;
       en        : in  std_logic;
       input     : in  std_logic_vector(wid-1 downto 0);
       output    : out std_logic_vector(wid-1 downto 0));
end REG;

architecture bhv of REG is
begin
  process(clk, rst)
  begin
    if rst = '1' then
      output   <= (others => init);
    elsif (clk = '1' and clk'event) then
      if (en = '1') then
        output <= input;
      end if;
    end if;
  end process;
end bhv;
