	 
	--******************************************************************************************
	--*  COMPANY    :  CHREC                                                                   *
	--*  NAME       :  Krishna Parthaje                                                        *
	--*  BOARD      :  PROCStarIV_530_1                                                        *
	--*  IC#        :  1                                                                       *
	--*  Created    :  Mon May 19 11:20:47 2014                                                *
	--*  This file  was  generated by  ProcWizard Application  version 9, 1, 2, 0              *
	--*  Copyright (C) 2014. All Rights Reserved to GiDEL Ltd                                  *
	--******************************************************************************************
	 
	 
	 
	 
	 
	 
	 
	 
	--======================================================================
	--=                   Use Altera Libraries For VHDL                    =
	--======================================================================
	LIBRARY altera;
	USE altera.altera_primitives_components.all;
	 
	 
	LIBRARY   ieee;
	USE       ieee.std_logic_1164.all;
	USE       ieee.std_logic_unsigned.all;
	USE       ieee.std_logic_arith.all;
	 
	ENTITY   tile   IS
	    PORT(

	--======================================================================
	--=                              Clocks                                =
	--======================================================================
		clk0                           : IN    STD_LOGIC;                          -- fast global clock
		clk2                           : IN    STD_LOGIC;                          -- slower global clock
		mem_ref_clk0                   : IN    STD_LOGIC;                          -- memory reference clock
		mem_ref_clk1                   : IN    STD_LOGIC;                          -- memory reference clock
	 
	--======================================================================
	--=                       Local Bus Connections                        =
	--======================================================================
		lb_rx                          : IN    STD_LOGIC_VECTOR( 32 DOWNTO 0 );    -- local bus data recieve
		lb_rx_clk                      : IN    STD_LOGIC;                          -- local bus recieve clock
		lb_tx                          : OUT   STD_LOGIC_VECTOR( 32 DOWNTO 0 );    -- local bus data transmit
		lb_tx_clk                      : OUT   STD_LOGIC;                          -- local bus transmit clock
		clrn                           : IN    STD_LOGIC;                          -- Device Global Clear Signal (active low)
		scl                            : IN    STD_LOGIC;                          -- Reserved I2C connection , do not use
		sda                            : IN    STD_LOGIC;                          -- Reserved I2C connection , do not use
	 
	--======================================================================
	--=                   DDR2 SDRAM block 1 (Onboard)                     =
	--======================================================================
		addr_a                         : OUT   STD_LOGIC_VECTOR( 13 DOWNTO 0 );    -- address bus
		ba_a                           : OUT   STD_LOGIC_VECTOR( 2  DOWNTO 0 );    -- bank address
		cas_a                          : OUT   STD_LOGIC;                          -- command input - active low
		cke_a                          : OUT   STD_LOGIC;                          -- clock enable  - active high
		ck_a                           : INOUT STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- clock
		ckn_a                          : INOUT STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- negative clock
		cs_a                           : OUT   STD_LOGIC;                          -- chip select   - active low
		dq_a                           : INOUT STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- data bus
		dqm_a                          : OUT   STD_LOGIC_VECTOR( 3  DOWNTO 0 );    -- output mask (byte enable)
		dqs_a                          : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- data strobe
		we_a                           : OUT   STD_LOGIC;                          -- command input - active low
		ras_a                          : OUT   STD_LOGIC;                          -- command input - active low
	 
	--======================================================================
	--=                    DDR2 SDRAM block 2 (SODIMM)                     =
	--======================================================================
		addr_b                         : OUT   STD_LOGIC_VECTOR( 15 DOWNTO 0 );    -- address bus
		ba_b                           : OUT   STD_LOGIC_VECTOR( 2  DOWNTO 0 );    -- bank address
		cas_b                          : OUT   STD_LOGIC;                          -- command input - active low
		cke_b                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- clock enable  - active high
		ck_b                           : INOUT STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- clock
		ckn_b                          : INOUT STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- negative clock
		cs_b                           : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- chip select   - active low
		dq_b                           : INOUT STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- data bus
		dqm_b                          : OUT   STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- output mask (byte enable)
		dqs_b                          : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- data strobe
		dqsn_b                         : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- negative data strobe
		we_b                           : OUT   STD_LOGIC;                          -- command input - active low
		ras_b                          : OUT   STD_LOGIC;                          -- command input - active low
		odt_b                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- built_in memory termination enable - active high
	 
	--======================================================================
	--=                    DDR2 SDRAM block 3 (SODIMM)                     =
	--======================================================================
		addr_c                         : OUT   STD_LOGIC_VECTOR( 15 DOWNTO 0 );    -- address bus
		ba_c                           : OUT   STD_LOGIC_VECTOR( 2  DOWNTO 0 );    -- bank address
		cas_c                          : OUT   STD_LOGIC;                          -- command input - active low
		cke_c                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- clock enable  - active high
		ck_c                           : INOUT STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- clock
		ckn_c                          : INOUT STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- negative clock
		cs_c                           : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- chip select   - active low
		dq_c                           : INOUT STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- data bus
		dqm_c                          : OUT   STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- output mask (byte enable)
		dqs_c                          : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- data strobe
		dqsn_c                         : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- negative data strobe
		we_c                           : OUT   STD_LOGIC;                          -- command input - active low
		ras_c                          : OUT   STD_LOGIC;                          -- command input - active low
		odt_c                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- built_in memory termination enable - active high
	 
	--======================================================================
	--=                       User Buses / Signals                         =
	--======================================================================
		v18_l                          : INOUT STD_LOGIC_VECTOR( 9  DOWNTO 0 );    -- 1.8V left bus
		v18_r                          : INOUT STD_LOGIC_VECTOR( 9  DOWNTO 0 );    -- 1.8V right bus
		main                           : INOUT STD_LOGIC_VECTOR( 39 DOWNTO 0 );    -- Common bus for IC1-IC4, MAIN(38:39) connected to J8,J10,J12,J14
		l                              : INOUT STD_LOGIC_VECTOR( 99 DOWNTO 0 );    -- Left bus
		l_in                           : IN    STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Left input bus connects to L connector
		l_io                           : INOUT STD_LOGIC_VECTOR( 19 DOWNTO 0 );    -- Left io bus connects to L connector
		clk_out                        : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock output to Left connector
		l2_l                           : INOUT STD_LOGIC_VECTOR( 84 DOWNTO 0 );    -- Second Left bus  connects to J12
		l2_in                          : IN    STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Second Left input bus  connects to J12
		l2_io                          : INOUT STD_LOGIC_VECTOR( 19 DOWNTO 0 );    -- Second Left io bus  connects to J12
		l2_clk_out                     : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Second clock output connects to J12
		led                            : OUT   STD_LOGIC_VECTOR( 3  DOWNTO 0 )     -- set '1' to light
	    );
	END   tile;
	 
	 
	ARCHITECTURE  tile_arch  OF  tile  IS
	CONSTANT    RBF_VERSION_VAL                       :STD_LOGIC_VECTOR := "00000001";
	 
	COMPONENT   tile_if
	    PORT(

	 
	--Local Bus Interface Signals
		clrn                           : IN    STD_LOGIC;                          -- User Global Clear   (0: clear all)
		lclk                           : OUT   STD_LOGIC;                          -- Local Bus Clock
		lb_rx_clk                      : IN    STD_LOGIC;                          -- Receiver (in) Local Bus Clock
		lb_rx                          : IN    STD_LOGIC_VECTOR( 32 DOWNTO 0 );    -- Local address/data bus (in)
		lb_tx_clk                      : OUT   STD_LOGIC;                          -- Transmitter (out) Local Bus Clock
		lb_tx                          : OUT   STD_LOGIC_VECTOR( 32 DOWNTO 0 );    -- Local address/data bus (out)
		g_reserved_control             : OUT   STD_LOGIC_VECTOR( 99 DOWNTO 0 );    -- Gidel reserved control bus (out)
		id                             : OUT   STD_LOGIC_VECTOR( 2  DOWNTO 0 );    -- FPGA number identification
	 
	--Internal Bus Interface Signals
		l_wr                           : OUT   STD_LOGIC;                          -- User Write Signal (1:write)
		addr_wr                        : OUT   STD_LOGIC_VECTOR( 31 DOWNTO 0 );    -- local bus address for write operations (including burst auto address increment)
		l_data_wr                      : OUT   STD_LOGIC_VECTOR( 127 DOWNTO 0 );   -- user input local data bus
		mem_ready_wr                   : IN    STD_LOGIC;                          -- 1: end of data write transfer (memory data is valid) on rising edge of lclk
		l_rd                           : OUT   STD_LOGIC;                          -- User Read Signal (0:read)
		addr_rd                        : OUT   STD_LOGIC_VECTOR( 31 DOWNTO 0 );    -- local bus address for read operations (including burst auto address increment)
		l_data_rd                      : IN    STD_LOGIC_VECTOR( 127 DOWNTO 0 );   -- data to read back from device memories
		mem_ready_rd                   : IN    STD_LOGIC;                          -- 1: end of data read transfer (memory data is valid) on rising edge of lclk
	 
	--Interrupt Logic
		interrupt                      : IN    STD_LOGIC;                          -- User interrupt
		interrupt_ack                  : OUT   STD_LOGIC;                          -- User interrupt acknowledge
	 
	--DREQ Logic
		user_dreq                      : IN    STD_LOGIC_VECTOR( 31 DOWNTO 0 );    -- User DMA control for each DMA channel
		done                           : IN    STD_LOGIC;
	 
	--version of RBF
		rbf_version                    : IN    STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- RBF_Info[7..0]
		almost_full_dst                : IN    STD_LOGIC;                          -- status_dst[1]
		go                             : OUT   STD_LOGIC;
		sel_reset_fifo                 : OUT   STD_LOGIC;                          -- select for reset_fifo
		sel_fifo_dst                   : OUT   STD_LOGIC;                          -- select for fifo_dst
		g_dreq_rd                      : IN    STD_LOGIC                           -- GiDEL DREQ signals
	    );
	END   COMPONENT;
	 
	 
	COMPONENT   user
	    PORT(

	 
	--Internal Bus Connections
		clrn                           : IN    STD_LOGIC;                          -- 0: global reset 
		clk0                           : IN    STD_LOGIC;                          -- Clock
		go                             : IN    STD_LOGIC;
		done                           : OUT   STD_LOGIC;
		Bank_A_ready                   : IN    STD_LOGIC;                          -- 1: Memory controller is ready for use, 0: Initializing (due to reset)
		data_src                       : OUT   STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- Data to the port src of FIFO fifo
		wr_req_fifo                    : OUT   STD_LOGIC;                          -- FIFO fifo write request signal
		wr_ack_fifo                    : IN    STD_LOGIC;                          -- FIFO fifo write acknowledge signal
		fifo_eos                       : IN    STD_LOGIC;                          -- 1: fifo port End of Stream pulse
		fifo_flush                     : OUT   STD_LOGIC;                          -- Flush FIFO data (assert high when the transfer is over)
		fifo_rewind                    : OUT   STD_LOGIC                           -- 1: Start read port from the beginning of the FIFO
	    );
	END   COMPONENT;
	 
	 
	COMPONENT   user_pll1
	    PORT(

		inclk0                         : IN    STD_LOGIC;
		c0                             : OUT   STD_LOGIC 
	    );
	END   COMPONENT;
	 
	 
	COMPONENT   IC_1_Bank_A_Ctrl
	    PORT(

	 
	--Global MultiPort Connections
		clrn                           : IN    STD_LOGIC;                          -- MultiPort async global reset
		ref_clk                        : IN    STD_LOGIC;                          -- SDRAM clock
		g_reserved_control             : IN    STD_LOGIC_VECTOR( 99 DOWNTO 0 );    -- SDRAM Connection
		ready                          : OUT   STD_LOGIC;                          -- 1: Memory controller is ready for use, 0: Initializing (due to reset)
	 
	--SDRAM Connections
		data                           : INOUT STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- Memory data
		addr                           : OUT   STD_LOGIC_VECTOR( 12 DOWNTO 0 );    -- Memory address
		dqm                            : OUT   STD_LOGIC_VECTOR( 3  DOWNTO 0 );    -- DQM signal from MultiPort
		dqs                            : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- DQS signal from MultiPort
		ba                             : OUT   STD_LOGIC_VECTOR( 2  DOWNTO 0 );    -- SDRAM control signal
		cs                             : OUT   STD_LOGIC;                          -- Chip Select signal from MultiPort 6
		ce                             : OUT   STD_LOGIC;                          -- Clock Enable signal from MultiPort 6
		ras                            : OUT   STD_LOGIC;                          -- RAS signal from MultiPort
		cas                            : OUT   STD_LOGIC;                          -- CAS signal from MultiPort
		we                             : OUT   STD_LOGIC;                          -- Write Enable signal from MultiPort
		ck                             : INOUT STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- CK
		ckn                            : INOUT STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- CKN
	 
	--Port src of FIFO fifo Connections
		clk_src                        : IN    STD_LOGIC;                          -- Port clock
		data_src                       : IN    STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- Data to the port src of FIFO fifo
		fifo_flush                     : IN    STD_LOGIC;                          -- Flush FIFO data (assert high when the transfer is over)
	 
	--Port dst of FIFO fifo Connections
		clk_dst                        : IN    STD_LOGIC;                          -- Port clock
		data_dst                       : OUT   STD_LOGIC_VECTOR( 127 DOWNTO 0 );   -- Data from the port dst of FIFO fifo
		fifo_almost_full_dst           : OUT   STD_LOGIC;                          -- MultiPort status to Host
	 
	--FIFO fifo Connections
		reset_fifo                     : IN    STD_LOGIC;                          -- FIFO fifo reset signal
		lclk                           : IN    STD_LOGIC;                          -- FIFO fifo reset signal clock
		sel_fifo                       : IN    STD_LOGIC;                          -- FIFO fifo read request from PCI
		wr_req_fifo                    : IN    STD_LOGIC;                          -- FIFO fifo write request signal
		wr_ack_fifo                    : OUT   STD_LOGIC;                          -- FIFO fifo write acknowledge signal
		almost_full_fifo               : OUT   STD_LOGIC;                          -- FIFO fifo almost full signal
		almost_empty_fifo              : OUT   STD_LOGIC;                          -- FIFO fifo almost empty signal
		half_full_fifo                 : OUT   STD_LOGIC;                          -- FIFO fifo half full signal
		g_dreq_fifo                    : OUT   STD_LOGIC;                          -- DMA transfer hold request from FIFO fifo
		fifo_eos                       : OUT   STD_LOGIC;                          -- 1: fifo port End of Stream pulse
		fifo_rewind                    : IN    STD_LOGIC                           -- 1: Start read port from the beginning of the FIFO
	    );
	END   COMPONENT;
	 
	 
	 
	 
	 
	--Local bus interfaces
	 
	--Hardware status registers (FPGA->Host)
	SIGNAL   done                       : STD_LOGIC;
	SIGNAL   rbf_version                : STD_LOGIC_VECTOR( 7  DOWNTO 0 );     -- RBF_Info[7..0]
	SIGNAL   almost_full_dst            : STD_LOGIC;                           -- status_dst[1]
	 
	--Mode registers (Host->FPGA). Use to set hardware working modes
	SIGNAL   g_reserved_control         : STD_LOGIC_VECTOR( 99 DOWNTO 0 );     -- Gidel reserved control bus
	SIGNAL   id                         : STD_LOGIC_VECTOR( 2  DOWNTO 0 );     -- FPGA number identification
	SIGNAL   lclk                       : STD_LOGIC;                           -- Local Bus Clock
	SIGNAL   l_wr                       : STD_LOGIC;                           -- User Write Signal (1:write)
	SIGNAL   addr_wr                    : STD_LOGIC_VECTOR( 31 DOWNTO 0 );     -- local bus address for write operations
	SIGNAL   l_data_wr                  : STD_LOGIC_VECTOR( 127 DOWNTO 0 );    -- user input local data bus
	SIGNAL   mem_ready_wr               : STD_LOGIC;                           -- 1: write memory data is valid (memory is ready)
	SIGNAL   l_rd                       : STD_LOGIC;                           -- User Read Signal (0:read)
	SIGNAL   addr_rd                    : STD_LOGIC_VECTOR( 31 DOWNTO 0 );     -- local bus address for read operations
	SIGNAL   l_data_rd                  : STD_LOGIC_VECTOR( 127 DOWNTO 0 );    -- data to read back from device memories
	SIGNAL   mem_ready_rd               : STD_LOGIC;                           -- 1: end of data read transfer (memory data is valid)
	 
	--User interrupt signals
	SIGNAL   interrupt                  : STD_LOGIC;                           -- Interrupt signal - assert low to send interrupt to SoftWare, when interrupt_ack is high.
	SIGNAL   interrupt_ack              : STD_LOGIC;                           -- Interrupt acknowledge signal - asserted high to to enable user interrupt.
	 
	--User DREQ signals
	SIGNAL   user_dreq                  : STD_LOGIC_VECTOR( 31 DOWNTO 0 );     -- DMA control - assert low to enable DMA operation, high to stop DMA (for each DMA channel).
	 
	--Other signals
	SIGNAL   go                         : STD_LOGIC;
	SIGNAL   clk                        : STD_LOGIC;
	 
	--Select signals for user's memories / reggroups
	SIGNAL   sel_reset_fifo             : STD_LOGIC;                           -- select for reset_fifo
	SIGNAL   sel_fifo_dst               : STD_LOGIC;                           -- select for fifo_dst
	 
	--FIFO fifo
	SIGNAL   Bank_A_ready               : STD_LOGIC;                           -- 1: Memory controller is ready for use, 0: Initializing (due to reset)
	SIGNAL   data_src                   : STD_LOGIC_VECTOR( 63 DOWNTO 0 );     -- Data to the port src of FIFO fifo
	SIGNAL   fifo_flush                 : STD_LOGIC;                           -- Flush FIFO data (assert high when the transfer is over)
	SIGNAL   data_dst                   : STD_LOGIC_VECTOR( 127 DOWNTO 0 );    -- Data from the port dst of FIFO fifo
	SIGNAL   wr_req_fifo                : STD_LOGIC;                           -- FIFO fifo write request signal
	SIGNAL   wr_ack_fifo                : STD_LOGIC;                           -- FIFO fifo write acknowledge signal
	SIGNAL   almost_full_fifo           : STD_LOGIC;                           -- FIFO fifo almost full signal
	SIGNAL   almost_empty_fifo          : STD_LOGIC;                           -- FIFO fifo almost empty signal
	SIGNAL   half_full_fifo             : STD_LOGIC;                           -- FIFO fifo half full signal
	SIGNAL   g_dreq_fifo                : STD_LOGIC;                           -- DMA transfer hold request from FIFO fifo
	SIGNAL   fifo_eos                   : STD_LOGIC;                           -- 1: fifo port End of Stream pulse
	SIGNAL   fifo_rewind                : STD_LOGIC;                           -- 1: Start read port from the beginning of the FIFO
	 
	 
	BEGIN
		 
		 
		 
		 
		--======================================================================
		--=    The Interface entity connections (connections to the host)      =
		--======================================================================
		if_tile : tile_if
		PORT MAP  (
		 
		--Local Bus Interface Signals
		clrn                         =>  clrn,                                     -- IN        User Global Clear   (0: clear all)
		lclk                         =>  lclk,                                     -- OUT       Local Bus Clock
		lb_rx_clk                    =>  lb_rx_clk,                                -- IN        Receiver (in) Local Bus Clock
		lb_rx( 32 DOWNTO 0 )         =>  lb_rx( 32 DOWNTO 0 ),                     -- IN        Local address/data bus (in)
		lb_tx_clk                    =>  lb_tx_clk,                                -- OUT       Transmitter (out) Local Bus Clock
		lb_tx( 32 DOWNTO 0 )         =>  lb_tx( 32 DOWNTO 0 ),                     -- OUT       Local address/data bus (out)
		g_reserved_control( 99 DOWNTO 0 )  =>  g_reserved_control( 99 DOWNTO 0 ),  -- OUT       Gidel reserved control bus (out)
		id( 2  DOWNTO 0 )            =>  id( 2  DOWNTO 0 ),                        -- OUT       FPGA number identification
		 
		--Internal Bus Interface Signals
		l_wr                         =>  l_wr,                                     -- OUT       User Write Signal (1:write)
		addr_wr( 31 DOWNTO 0 )       =>  addr_wr( 31 DOWNTO 0 ),                   -- OUT       local bus address for write operations (including burst auto address increment)
		l_data_wr( 127 DOWNTO 0 )    =>  l_data_wr( 127 DOWNTO 0 ),                -- OUT       user input local data bus
		mem_ready_wr                 =>  mem_ready_wr,                             -- IN        1: end of data write transfer (memory data is valid) on rising edge of lclk
		l_rd                         =>  l_rd,                                     -- OUT       User Read Signal (0:read)
		addr_rd( 31 DOWNTO 0 )       =>  addr_rd( 31 DOWNTO 0 ),                   -- OUT       local bus address for read operations (including burst auto address increment)
		l_data_rd( 127 DOWNTO 0 )    =>  l_data_rd( 127 DOWNTO 0 ),                -- IN        data to read back from device memories
		mem_ready_rd                 =>  mem_ready_rd,                             -- IN        1: end of data read transfer (memory data is valid) on rising edge of lclk
		 
		--Interrupt Logic
		interrupt                    =>  interrupt,                                -- IN        User interrupt
		interrupt_ack                =>  interrupt_ack,                            -- OUT       User interrupt acknowledge
		 
		--DREQ Logic
		user_dreq( 31 DOWNTO 0 )     =>  user_dreq( 31 DOWNTO 0 ),                 -- IN        User DMA control for each DMA channel
		 
		--Hardware status registers (FPGA->Host)
		done                         =>  done,                                     -- IN   
		rbf_version( 7  DOWNTO 0 )   =>  rbf_version( 7  DOWNTO 0 ),               -- IN        RBF_Info[7..0]
		almost_full_dst              =>  almost_full_dst,                          -- IN        status_dst[1]
		 
		--Mode registers (Host->FPGA). Use to set hardware working modes
		go                           =>  go,                                       -- OUT  
		 
		--Select signals for user's memories / reggroups
		sel_reset_fifo               =>  sel_reset_fifo,                           -- OUT       select for reset_fifo
		sel_fifo_dst                 =>  sel_fifo_dst,                             -- OUT       select for fifo_dst
		g_dreq_rd                    =>  g_dreq_fifo                               -- IN   
		);

		 
		 
		 
		 
		--======================================================================
		--=                   User's entities' connections                     =
		--======================================================================
		 
		 
		--user
		 
		user_cmp : user
		PORT MAP  (
		clrn                         =>  clrn,                                     -- IN   
		clk0                         =>  clk0,                                     -- IN   
		go                           =>  go,                                       -- IN   
		done                         =>  done,                                     -- OUT  
		Bank_A_ready                 =>  Bank_A_ready,                             -- IN        1: Memory controller is ready for use, 0: Initializing (due to reset)
		data_src                     =>  data_src,                                 -- OUT       Data to the port src of FIFO fifo
		wr_req_fifo                  =>  wr_req_fifo,                              -- OUT       FIFO fifo write request signal
		wr_ack_fifo                  =>  wr_ack_fifo,                              -- IN        FIFO fifo write acknowledge signal
		fifo_eos                     =>  fifo_eos,                                 -- IN        1: fifo port End of Stream pulse
		fifo_flush                   =>  fifo_flush,                               -- OUT       Flush FIFO data (assert high when the transfer is over)
		fifo_rewind                  =>  fifo_rewind                               -- OUT       1: Start read port from the beginning of the FIFO
		);

		 
		 
		 
		--*********** FINISH *************
		 
		 
		 
		 
		--======================================================================
		--=                      User PLLs' connections                        =
		--======================================================================
		 
		user_pll1_cmp : user_pll1
		PORT MAP  (
		inclk0                       =>  clk0,                                     -- IN   
		c0                           =>  clk                                       -- OUT       250.000000 MHz @ 0.000000 deg.
		);

		 
		 
		 
		 
		--======================================================================
		--=                   SDRAM controllers' connections                   =
		--======================================================================
		 
		--======================================================================
		--=                         IC_1_Bank_A_Ctrl                           =
		--======================================================================
		 
		 
		IC_1_Bank_A_Ctrl_cmp : IC_1_Bank_A_Ctrl
		PORT MAP  (
		 
		--Global MultiPort Connections
		clrn                         =>  clrn,                                     -- IN   
		ref_clk                      =>  mem_ref_clk0,                             -- IN   
		g_reserved_control( 99 DOWNTO 0 )  =>  g_reserved_control( 99 DOWNTO 0 ),  -- IN   
		ready                        =>  Bank_A_ready,                             -- OUT  
		 
		--SDRAM Connections
		data( 63 DOWNTO 0 )          =>  dq_a( 63 DOWNTO 0 ),                      -- OUT  
		addr( 12 DOWNTO 0 )          =>  addr_a( 12 DOWNTO 0 ),                    -- OUT  
		dqm( 3  DOWNTO 0 )           =>  dqm_a( 3  DOWNTO 0 ),                     -- OUT  
		dqs( 7  DOWNTO 0 )           =>  dqs_a( 7  DOWNTO 0 ),                     -- OUT  
		ba( 2  DOWNTO 0 )            =>  ba_a( 2  DOWNTO 0 ),                      -- OUT  
		cs                           =>  cs_a,                                     -- OUT  
		ce                           =>  cke_a,                                    -- OUT  
		ras                          =>  ras_a,                                    -- OUT  
		cas                          =>  cas_a,                                    -- OUT  
		we                           =>  we_a,                                     -- OUT  
		ck( 1  DOWNTO 0 )            =>  ck_a( 1  DOWNTO 0 ),                      -- OUT  
		ckn( 1  DOWNTO 0 )           =>  ckn_a( 1  DOWNTO 0 ),                     -- OUT  
		 
		--Port src of FIFO fifo Connections
		clk_src                      =>  clk0,                                     -- IN   
		data_src( 63 DOWNTO 0 )      =>  data_src( 63 DOWNTO 0 ),                  -- IN   
		fifo_flush                   =>  fifo_flush,                               -- IN   
		 
		--Port dst of FIFO fifo Connections
		clk_dst                      =>  lclk,                                     -- IN   
		data_dst( 127 DOWNTO 0 )     =>  data_dst( 127 DOWNTO 0 ),                 -- OUT  
		fifo_almost_full_dst         =>  almost_full_dst,                          -- OUT  
		 
		--FIFO fifo Connections
		reset_fifo                   =>  sel_reset_fifo,                           -- IN   
		lclk                         =>  lclk,                                     -- IN   
		sel_fifo                     =>  sel_fifo_dst,                             -- IN   
		wr_req_fifo                  =>  wr_req_fifo,                              -- IN   
		wr_ack_fifo                  =>  wr_ack_fifo,                              -- OUT  
		almost_full_fifo             =>  almost_full_fifo,                         -- OUT  
		almost_empty_fifo            =>  almost_empty_fifo,                        -- OUT  
		half_full_fifo               =>  half_full_fifo,                           -- OUT  
		g_dreq_fifo                  =>  g_dreq_fifo,                              -- OUT  
		fifo_eos                     =>  fifo_eos,                                 -- OUT  
		fifo_rewind                  =>  fifo_rewind                               -- IN   
		);

		 
		 
		rbf_version(7 DOWNTO 0)    <=    RBF_VERSION_VAL;  
		 
		 
		--======================================================================
		--=                Default Values of Board Connections                 =
		--======================================================================
		 
		--DDR Block B Connections
		addr_b                       <=  ( others => '0' );
		ba_b                         <=  ( others => '0' );
		cas_b                        <=  '0';
		cke_b                        <=  ( others => '0' );
		ck_b                         <=  ( others => 'Z' );
		ckn_b                        <=  ( others => 'Z' );
		cs_b                         <=  ( others => '1' );
		dq_b                         <=  ( others => 'Z' );
		dqm_b                        <=  ( others => '0' );
		dqs_b                        <=  ( others => 'Z' );
		dqsn_b                       <=  ( others => 'Z' );
		we_b                         <=  '0';
		ras_b                        <=  '0';
		odt_b                        <=  ( others => '0' );
		 
		--DDR Block C Connections
		addr_c                       <=  ( others => '0' );
		ba_c                         <=  ( others => '0' );
		cas_c                        <=  '0';
		cke_c                        <=  ( others => '0' );
		ck_c                         <=  ( others => 'Z' );
		ckn_c                        <=  ( others => 'Z' );
		cs_c                         <=  ( others => '1' );
		dq_c                         <=  ( others => 'Z' );
		dqm_c                        <=  ( others => '0' );
		dqs_c                        <=  ( others => 'Z' );
		dqsn_c                       <=  ( others => 'Z' );
		we_c                         <=  '0';
		ras_c                        <=  '0';
		odt_c                        <=  ( others => '0' );
		 
		--User's buses
		 
		mem_ready_wr                 <=  '1';                                      -- '1'   NO WAIT STATES, put '0' when you want to add wait states
		 
		mem_ready_rd                 <=  '1';                                      -- '1'   NO WAIT STATES, put '0' when you want to add wait states
		l_data_rd( 31 DOWNTO 0 )     <= data_dst( 31 DOWNTO 0 )   ;
		 
		l_data_rd( 127 DOWNTO 32 )   <= data_dst( 127 DOWNTO 32 )   ;
		 
		interrupt                    <=  '1';                                      -- Interrupt control - assert low to send interrupt to SoftWare, when interrupt_ack is high.
		user_dreq                    <=  ( others => '0' );                        -- DMA control - assert low to enable DMA operation, high to stop DMA (for each DMA channel).
		v18_l                        <=  ( others => 'Z' );
		v18_r                        <=  ( others => 'Z' );
		main                         <=  ( others => 'Z' );
		l                            <=  ( others => 'Z' );
		l_io                         <=  ( others => 'Z' );
		clk_out                      <=  ( others => '0' );
		l2_l                         <=  ( others => 'Z' );
		l2_io                        <=  ( others => 'Z' );
		led                          <=  ( others => '0' );
		 
		 
	END  tile_arch;
