	 
	--******************************************************************************************
	--*  COMPANY    :  ________                                                                *
	--*  NAME       :  Krishna                                                                 *
	--*  BOARD      :  ProceV_D8                                                               *
	--*  IC#        :  1                                                                       *
	--*  Created    :  Fri Jan 23 09:27:18 2015                                                *
	--*  This file  was  generated by  ProcWizard Application  version 9.2.1.0                 *
	--*  Copyright (C) 2015. All Rights Reserved to GiDEL Ltd                                  *
	--******************************************************************************************
	 
	 
	 
	 
	 
	 
	 
	 
	--======================================================================
	--=                   Use Altera Libraries For VHDL                    =
	--======================================================================
	LIBRARY altera;
	USE altera.altera_primitives_components.all;
	 
	 
	LIBRARY   ieee;
	USE       ieee.std_logic_1164.all;
	USE       ieee.std_logic_unsigned.all;
	USE       ieee.std_logic_arith.all;
	 
	ENTITY   tile   IS
	    PORT(

	--======================================================================
	--=                         Clocks & Globals                           =
	--======================================================================
		ref_clk                        : IN    STD_LOGIC;                          -- 25 MHz reference clock input pin
		mem_ref_clk                    : IN    STD_LOGIC;                          -- 125MHz, memory reference clock input pin
		ext_clk                        : IN    STD_LOGIC;                          -- User external clock from SMA
		ext_resetn                     : IN    STD_LOGIC;                          -- Used in stand-alone from push button
		scl                            : INOUT STD_LOGIC;                          -- SODIMM Serial clock. Used to synchronize communication to and from the I2C bus
		sda                            : INOUT STD_LOGIC;                          -- SODIMM Serial data:  Used to transfer addresses and data into and out of the I2C bus
		ledn                           : OUT   STD_LOGIC_VECTOR( 4  DOWNTO 1 );    -- General Purpose User LEDs; 0: light on
		status_ledn                    : OUT   STD_LOGIC_VECTOR( 3  DOWNTO 1 );    -- Status LEDs; 0: light on
		g_reserved                     : INOUT STD_LOGIC_VECTOR( 33 DOWNTO 0 );    -- Gidel reserved IO bus
	 
	--======================================================================
	--=                       PCIe Bus Connections                         =
	--======================================================================
		pcie_refclk                    : IN    STD_LOGIC;                          -- Reference clock for the Stratix V Hard IP for PCI Express
		pcie_perst                     : IN    STD_LOGIC;                          -- Active low reset from the PCIe reset pin of the device
		pcie_rx                        : IN    STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Receive inputs. These signals are the serial inputs of lanes 7�0
		pcie_tx                        : OUT   STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Transmit outputs. These signals are the serial outputs of lanes 7�0
	 
	--======================================================================
	--=                    DDR3 SDRAM block B (SODIMM)                     =
	--======================================================================
		addr_b                         : OUT   STD_LOGIC_VECTOR( 15 DOWNTO 0 );    -- Address bus
		ba_b                           : OUT   STD_LOGIC_VECTOR( 2  DOWNTO 0 );    -- Bank address select
		cas_b                          : OUT   STD_LOGIC;                          -- Command output(CAS) - active LOW
		cke_b                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock enable - active HIGH
		ck_b                           : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock: Differential clock outputs (positive)
		ckn_b                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock: Differential clock outputs (negative)
		cs_b                           : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Chip select - active LOW
		dq_b                           : INOUT STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- Data bus
		dqm_b                          : OUT   STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Data mask,is an output mask signal for write data (byte enable)
		dqs_b                          : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Data strobe: Differential data strobes (positive)
		dqsn_b                         : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Data strobe: Differential data strobes (negative)
		we_b                           : OUT   STD_LOGIC;                          -- Write enable - active LOW
		ras_b                          : OUT   STD_LOGIC;                          -- Command output(RAS) - active LOW
		odt_b                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- On-die termination enable - active HIGH
		resetn_b                       : OUT   STD_LOGIC;                          -- asynchronous SODIMM Reset - active LOW
		event_b                        : IN    STD_LOGIC;                          -- 1: SODIMM critical temperature thresholds have been exceeded
		rzq_b                          : IN    STD_LOGIC;                          -- Used for OCT calibration, the RZQ pin is connected to GND through an external 240-Ohm reference resistor
	 
	--======================================================================
	--=                    DDR3 SDRAM block C (SODIMM)                     =
	--======================================================================
		addr_c                         : OUT   STD_LOGIC_VECTOR( 15 DOWNTO 0 );    -- Address bus
		ba_c                           : OUT   STD_LOGIC_VECTOR( 2  DOWNTO 0 );    -- Bank address select
		cas_c                          : OUT   STD_LOGIC;                          -- Command output(CAS) - active LOW
		cke_c                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock enable - active HIGH
		ck_c                           : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock: Differential clock outputs (positive)
		ckn_c                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock: Differential clock outputs (negative)
		cs_c                           : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Chip select - active LOW
		dq_c                           : INOUT STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- Data bus
		dqm_c                          : OUT   STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Data mask,is an output mask signal for write data (byte enable)
		dqs_c                          : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Data strobe: Differential data strobes (positive)
		dqsn_c                         : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Data strobe: Differential data strobes (negative)
		we_c                           : OUT   STD_LOGIC;                          -- Write enable - active LOW
		ras_c                          : OUT   STD_LOGIC;                          -- Command output(RAS) - active LOW
		odt_c                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- On-die termination enable - active HIGH
		resetn_c                       : OUT   STD_LOGIC;                          -- asynchronous SODIMM Reset - active LOW
		event_c                        : IN    STD_LOGIC;                          -- 1: SODIMM critical temperature thresholds have been exceeded
		rzq_c                          : IN    STD_LOGIC;                          -- Used for OCT calibration, the RZQ pin is connected to GND through an external 240-Ohm reference resistor
	 
	--======================================================================
	--=                    DDR2 SRAM block D (Onboard)                     =
	--======================================================================
		dq_d                           : INOUT STD_LOGIC_VECTOR( 35 DOWNTO 0 );    -- Data bus
		ldn_d                          : OUT   STD_LOGIC;                          -- Synchronous load - active LOW
		bwsn_d                         : OUT   STD_LOGIC_VECTOR( 3  DOWNTO 0 );    -- Byte Write Select - active LOW
		r_wn_d                         : OUT   STD_LOGIC;                          -- 1: Synchronous read 0: Synchronous write
		k_d                            : OUT   STD_LOGIC;                          -- Positive output clock input
		cq_d                           : IN    STD_LOGIC;                          -- Clock (positive) synchronized to the input data
		cqn_d                          : IN    STD_LOGIC;                          -- Do not use
		qvld_d                         : IN    STD_LOGIC;                          -- 1: valid input data. QVLD is edge aligned with CQ and CQn.
		addr_d                         : OUT   STD_LOGIC_VECTOR( 21 DOWNTO 0 );    -- Address bus
	 
	--======================================================================
	--=                    DDR2 SRAM block E (Onboard)                     =
	--======================================================================
		dq_e                           : INOUT STD_LOGIC_VECTOR( 35 DOWNTO 0 );    -- Data bus
		ldn_e                          : OUT   STD_LOGIC;                          -- Synchronous load - active LOW
		bwsn_e                         : OUT   STD_LOGIC_VECTOR( 3  DOWNTO 0 );    -- Byte Write Select - active LOW
		r_wn_e                         : OUT   STD_LOGIC;                          -- 1: Synchronous read 0: Synchronous write
		k_e                            : OUT   STD_LOGIC;                          -- Positive output clock input
		cq_e                           : IN    STD_LOGIC;                          -- Clock (positive) synchronized to the input data
		cqn_e                          : IN    STD_LOGIC;                          -- Do not use
		qvld_e                         : IN    STD_LOGIC;                          -- 1: valid input data. QVLD is edge aligned with CQ and CQn.
		addr_e                         : OUT   STD_LOGIC_VECTOR( 21 DOWNTO 0 );    -- Address bus
	 
	--======================================================================
	--=                       User Buses / Signals                         =
	--======================================================================
	--======================================================================
	--=            1G PHY I/O's (Connections to on board PHY)              =
	--======================================================================
		phy_mdio                       : INOUT STD_LOGIC;                          -- Is a management data
		phy_mdc                        : OUT   STD_LOGIC;                          -- Is a management data clock reference
		phy_resetn                     : OUT   STD_LOGIC;                          -- Is a hardware reset - active LOW
		phy_rx_ctrl                    : IN    STD_LOGIC;                          -- Is a RGMII receive control
		phy_rx_clk                     : IN    STD_LOGIC;                          -- Is a RGMII receive clock
		phy_rxd                        : IN    STD_LOGIC_VECTOR( 3  DOWNTO 0 );    -- Is a RGMII receive data
		phy_tx_ctrl                    : OUT   STD_LOGIC;                          -- Is a RGMII transmit control
		phy_tx_clk                     : OUT   STD_LOGIC;                          -- Is a RGMII transmit clock
		phy_txd                        : OUT   STD_LOGIC_VECTOR( 3  DOWNTO 0 );    -- Is a RGMII transmit data
	 
	--======================================================================
	--=                               SFP A                                =
	--======================================================================
		sfp_mod_abs_a                  : IN    STD_LOGIC;                          -- 0: Module Absent, 1: Module inserted
		sfp_link_ledn_a                : OUT   STD_LOGIC;                          -- 0: led on
		sfp_trafic_ledn_a              : OUT   STD_LOGIC;                          -- 0: led on
	--======================================================================
	--=                               SFP B                                =
	--======================================================================
		sfp_mod_abs_b                  : IN    STD_LOGIC;                          -- 0: Module Absent, 1: Module inserted
		sfp_link_ledn_b                : OUT   STD_LOGIC;                          -- 0: led on
		sfp_trafic_ledn_b              : OUT   STD_LOGIC;                          -- 0: led on
	 
	--======================================================================
	--=                                CXP                                 =
	--======================================================================
		cxp_prsnt_l                    : IN    STD_LOGIC;                          -- Is used to indicate when the module is plugged into the host receptacle
	--======================================================================
	--=       High Speed (HS-B) - 8 lanes transceivers connections         =
	--======================================================================
		hs_prsnt_b                     : IN    STD_LOGIC;                          -- 0: This port is connected
	--======================================================================
	--=       High Speed (HS-C) - 4 lanes transceivers connections         =
	--======================================================================
		hs_prsnt_c                     : IN    STD_LOGIC;                          -- 0: This port is connected
	--======================================================================
	--=                   External(J3) connector I/O's                     =
	--======================================================================
		j3_ext_io                      : INOUT STD_LOGIC_VECTOR( 11 DOWNTO 0 );    -- General-purpose I/O bus
		j3_ext_io_dir                  : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Bit-0 sets direction for ext_io[7:0] and bit-1 for ext_io[11:8]. (ext_io_dir=0: Inputs, ext_io_dir=1: Outputs)
	--======================================================================
	--=                       L(J4) connector I/O's                        =
	--======================================================================
		l                              : INOUT STD_LOGIC_VECTOR( 84 DOWNTO 0 );    -- Bidirectional Left bus
		l_in                           : IN    STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Left input bus
		l_io                           : INOUT STD_LOGIC_VECTOR( 19 DOWNTO 0 );    -- Left io bus
		clk_out                        : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 )     -- Clock output
	    );
	END   tile;
	 
	 
	ARCHITECTURE  tile_arch  OF  tile  IS
	CONSTANT    RBF_VERSION_VAL                       :STD_LOGIC_VECTOR := "00000001";
	 
	COMPONENT   tile_if
	    PORT(

	 
	--Clocks & Globals
		ref_clk                        : IN    STD_LOGIC;                          -- 25 MHz reference clock input pin
		clk0                           : OUT   STD_LOGIC;                          -- Main system clock, the max frequency is 300 MHZ
		clk                            : OUT   STD_LOGIC;                          -- User clock, the frequency is twice/triply the frequency of clk0
		clk2                           : OUT   STD_LOGIC;                          -- Is an auxiliary clock that may be used as a slow emulation clock
		mem_ref_clk_int                : OUT   STD_LOGIC;                          -- Is an internal (from PLL) memory reference clock (125MHz)
		scl                            : INOUT STD_LOGIC;                          -- Serial clock. Used to synchronize communication to and from the I2C bus
		sda                            : INOUT STD_LOGIC;                          -- Serial data: Used to transfer addresses and data into and out of the I2C bus
		status_ledn                    : OUT   STD_LOGIC_VECTOR( 3  DOWNTO 1 );    -- Status LEDs; 0: light on
		id                             : OUT   STD_LOGIC_VECTOR( 2  DOWNTO 0 );    -- FPGA number identification
		g_reserved                     : INOUT STD_LOGIC_VECTOR( 33 DOWNTO 0 );    -- Gidel reserved IO bus
		g_reserved_control             : OUT   STD_LOGIC_VECTOR( 99 DOWNTO 0 );    -- Gidel reserved control bus (out)
	 
	--PCIe connection
		pcie_refclk                    : IN    STD_LOGIC;                          -- Reference clock for the Hard IP for PCI Express
		pcie_perst                     : IN    STD_LOGIC;                          -- Active low reset from the PCIe reset pin of the device
		pcie_rx                        : IN    STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Receive inputs. These signals are the serial inputs of lanes 7�0
		pcie_tx                        : OUT   STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Transmit outputs. These signals are the serial outputs of lanes 7�0
	 
	--Internal Bus Interface Signals
		clrn                           : OUT   STD_LOGIC;                          -- User Global Clear   (0: clear all)
		lclk                           : OUT   STD_LOGIC;                          -- Local Bus Clock
		l_wr                           : OUT   STD_LOGIC;                          -- User Write Signal (1:write)
		addr_wr                        : OUT   STD_LOGIC_VECTOR( 31 DOWNTO 0 );    -- local bus address for write operations (including burst auto address increment)
		l_data_wr                      : OUT   STD_LOGIC_VECTOR( 255 DOWNTO 0 );   -- user input local data bus
		mem_ready_wr                   : IN    STD_LOGIC;                          -- 1: end of data write transfer (memory data is valid) on rising edge of lclk
		l_rd                           : OUT   STD_LOGIC;                          -- User Read Signal (0:read)
		addr_rd                        : OUT   STD_LOGIC_VECTOR( 31 DOWNTO 0 );    -- local bus address for read operations (including burst auto address increment)
		l_data_rd                      : IN    STD_LOGIC_VECTOR( 255 DOWNTO 0 );   -- data to read back from device memories
		mem_ready_rd                   : IN    STD_LOGIC;                          -- 1: end of data read transfer (memory data is valid) on rising edge of lclk
	 
	--Interrupt Logic
		interrupt                      : IN    STD_LOGIC;                          -- User interrupt
		interrupt_ack                  : OUT   STD_LOGIC;                          -- User interrupt acknowledge
	 
	--DREQ Logic
		user_dreq                      : IN    STD_LOGIC_VECTOR( 31 DOWNTO 0 );    -- User DMA control for each DMA channel
		done                           : IN    STD_LOGIC;
	 
	--version of RBF
		rbf_version                    : IN    STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- RBF_Info[7..0]
		almost_full_dst                : IN    STD_LOGIC;                          -- status_dst[1]
		go                             : OUT   STD_LOGIC;
		sel_reset_singlea              : OUT   STD_LOGIC;                          -- select for reset_singlea
		sel_singlea_dst                : OUT   STD_LOGIC;                          -- select for singlea_dst
		g_dreq_rd                      : IN    STD_LOGIC                           -- GiDEL DREQ signals
	    );
	END   COMPONENT;
	 
	 
	 
	--g_mp_pll_sv
	COMPONENT   g_mp_pll_sv
	    PORT(

		clrn                           : IN    STD_LOGIC;
		mem_ref_clk                    : IN    STD_LOGIC;
		pll_mem_clk                    : OUT   STD_LOGIC;
		pll_write_clk                  : OUT   STD_LOGIC;
		pll_write_clk_pre_phy_clk      : OUT   STD_LOGIC;
		pll_addr_cmd_clk               : OUT   STD_LOGIC;
		pll_hr_clk                     : OUT   STD_LOGIC;
		pll_p2c_read_clk               : OUT   STD_LOGIC;
		pll_c2p_write_clk              : OUT   STD_LOGIC;
		pll_avl_clk                    : OUT   STD_LOGIC;
		pll_config_clk                 : OUT   STD_LOGIC;
		pll_locked                     : OUT   STD_LOGIC;
		afi_clk                        : OUT   STD_LOGIC;
		afi_half_clk                   : OUT   STD_LOGIC 
	    );
	END   COMPONENT;
	 
	 
	 
	 
	COMPONENT   user
	    PORT(

	 
	--Internal Bus Connections
		clrn                           : IN    STD_LOGIC;                          -- 0: global reset 
		clk0                           : IN    STD_LOGIC;                          -- Clock
		go                             : IN    STD_LOGIC;
		done                           : OUT   STD_LOGIC;
		Bank_B_ready                   : IN    STD_LOGIC;                          -- 1: Memory controller is ready for use, 0: Initializing (due to reset)
		data_src                       : OUT   STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- Data to the port src of FIFO singlea
		wr_req_singlea                 : OUT   STD_LOGIC;                          -- FIFO singlea write request signal
		wr_ack_singlea                 : IN    STD_LOGIC;                          -- FIFO singlea write acknowledge signal
		singlea_eos                    : IN    STD_LOGIC;                          -- 1: singlea port End of Stream pulse
		singlea_flush                  : OUT   STD_LOGIC;                          -- Flush FIFO data (assert high when the transfer is over)
		singlea_rewind                 : OUT   STD_LOGIC                           -- 1: Start read port from the beginning of the FIFO
	    );
	END   COMPONENT;
	 
	 
	COMPONENT   IC_1_Bank_B_Ctrl
	    PORT(

	 
	--Global MultiPort Connections
		clrn                           : IN    STD_LOGIC;                          -- MultiPort async global reset
		ref_clk                        : IN    STD_LOGIC;                          -- mem ref clock
		pll_mem_clk                    : IN    STD_LOGIC;
		pll_write_clk                  : IN    STD_LOGIC;
		pll_write_clk_pre_phy_clk      : IN    STD_LOGIC;
		pll_addr_cmd_clk               : IN    STD_LOGIC;
		pll_hr_clk                     : IN    STD_LOGIC;
		pll_p2c_read_clk               : IN    STD_LOGIC;
		pll_c2p_write_clk              : IN    STD_LOGIC;
		pll_avl_clk                    : IN    STD_LOGIC;
		pll_config_clk                 : IN    STD_LOGIC;
		pll_locked                     : IN    STD_LOGIC;
		afi_clk                        : IN    STD_LOGIC;
		afi_half_clk                   : IN    STD_LOGIC;
		g_reserved_control             : IN    STD_LOGIC_VECTOR( 99 DOWNTO 0 );    -- SDRAM Connection
		ready                          : OUT   STD_LOGIC;                          -- 1: Memory controller is ready for use, 0: Initializing (due to reset)
	 
	--SDRAM Connections
		data                           : INOUT STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- Memory data
		addr                           : OUT   STD_LOGIC_VECTOR( 15 DOWNTO 0 );    -- Memory address
		dqm                            : OUT   STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- DQM signal from MultiPort
		dqs                            : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- DQS signal from MultiPort
		dqsn                           : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- DQSN signal from MultiPort
		ba                             : OUT   STD_LOGIC_VECTOR( 2  DOWNTO 0 );    -- SDRAM control signal
		cs_bus                         : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Chip Select signal from MultiPort 4
		ce                             : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock Enable signal from MultiPort
		ras                            : OUT   STD_LOGIC;                          -- RAS signal from MultiPort
		cas                            : OUT   STD_LOGIC;                          -- CAS signal from MultiPort
		we                             : OUT   STD_LOGIC;                          -- Write Enable signal from MultiPort
		odt                            : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- ODT signal from MultiPort
		ck                             : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- CK
		ckn                            : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- CKN
		oct_rzqin                      : IN    STD_LOGIC;                          -- RZK signal from MultiPort
		event_in                       : IN    STD_LOGIC;                          -- event signal from MultiPort
		mem_reset_n                    : OUT   STD_LOGIC;                          -- resetn signal from MultiPort
	 
	--Port src of FIFO singlea Connections
		clk_src                        : IN    STD_LOGIC;                          -- Port clock
		data_src                       : IN    STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- Data to the port src of FIFO singlea
		singlea_flush                  : IN    STD_LOGIC;                          -- Flush FIFO data (assert high when the transfer is over)
	 
	--Port dst of FIFO singlea Connections
		clk_dst                        : IN    STD_LOGIC;                          -- Port clock
		data_dst                       : OUT   STD_LOGIC_VECTOR( 255 DOWNTO 0 );   -- Data from the port dst of FIFO singlea
		singlea_almost_full_dst        : OUT   STD_LOGIC;                          -- MultiPort status to Host
	 
	--FIFO singlea Connections
		reset_singlea                  : IN    STD_LOGIC;                          -- FIFO singlea reset signal
		lclk                           : IN    STD_LOGIC;                          -- FIFO singlea reset signal clock
		sel_singlea                    : IN    STD_LOGIC;                          -- FIFO singlea read request from PCI
		wr_req_singlea                 : IN    STD_LOGIC;                          -- FIFO singlea write request signal
		wr_ack_singlea                 : OUT   STD_LOGIC;                          -- FIFO singlea write acknowledge signal
		almost_full_singlea            : OUT   STD_LOGIC;                          -- FIFO singlea almost full signal
		almost_empty_singlea           : OUT   STD_LOGIC;                          -- FIFO singlea almost empty signal
		half_full_singlea              : OUT   STD_LOGIC;                          -- FIFO singlea half full signal
		g_dreq_singlea                 : OUT   STD_LOGIC;                          -- DMA transfer hold request from FIFO singlea
		singlea_eos                    : OUT   STD_LOGIC;                          -- 1: singlea port End of Stream pulse
		singlea_rewind                 : IN    STD_LOGIC                           -- 1: Start read port from the beginning of the FIFO
	    );
	END   COMPONENT;
	 
	 
	 
	 
	--Clocks & Globals
	 
	--Hardware status registers (FPGA->Host)
	SIGNAL   done                       : STD_LOGIC;
	SIGNAL   rbf_version                : STD_LOGIC_VECTOR( 7  DOWNTO 0 );     -- RBF_Info[7..0]
	SIGNAL   almost_full_dst            : STD_LOGIC;                           -- status_dst[1]
	 
	--Mode registers (Host->FPGA). Use to set hardware working modes
	SIGNAL   clk0                       : STD_LOGIC;                           -- Main system clock, the max frequency is 300 MHZ
	SIGNAL   clk                        : STD_LOGIC;                           -- User clock, the frequency is twice/triply the frequency of clk0
	SIGNAL   clk2                       : STD_LOGIC;                           -- Is an auxiliary clock that may be used as a slow emulation clock
	SIGNAL   mem_ref_clk_int            : STD_LOGIC;                           -- Is an internal (from PLL) memory reference clock (125MHz)
	SIGNAL   id                         : STD_LOGIC_VECTOR( 2  DOWNTO 0 );     -- FPGA number identification
	SIGNAL   g_reserved_control         : STD_LOGIC_VECTOR( 99 DOWNTO 0 );     -- Gidel reserved control bus
	 
	--Internal Bus Interface Signals
	SIGNAL   clrn                       : STD_LOGIC;                           -- User Global Clear   (0: clear all)
	SIGNAL   lclk                       : STD_LOGIC;                           -- Local Bus Clock
	SIGNAL   l_wr                       : STD_LOGIC;                           -- User Write Signal (1:write)
	SIGNAL   addr_wr                    : STD_LOGIC_VECTOR( 31 DOWNTO 0 );     -- local bus address for write operations
	SIGNAL   l_data_wr                  : STD_LOGIC_VECTOR( 255 DOWNTO 0 );    -- user input local data bus
	SIGNAL   mem_ready_wr               : STD_LOGIC;                           -- 1: write memory data is valid (memory is ready)
	SIGNAL   l_rd                       : STD_LOGIC;                           -- User Read Signal (0:read)
	SIGNAL   addr_rd                    : STD_LOGIC_VECTOR( 31 DOWNTO 0 );     -- local bus address for read operations
	SIGNAL   l_data_rd                  : STD_LOGIC_VECTOR( 255 DOWNTO 0 );    -- data to read back from device memories
	SIGNAL   mem_ready_rd               : STD_LOGIC;                           -- 1: end of data read transfer (memory data is valid)
	 
	--User interrupt signals
	SIGNAL   interrupt                  : STD_LOGIC;                           -- Interrupt signal - assert low to send interrupt to SoftWare, when interrupt_ack is high.
	SIGNAL   interrupt_ack              : STD_LOGIC;                           -- Interrupt acknowledge signal - asserted high to to enable user interrupt.
	 
	--User DREQ signals
	SIGNAL   user_dreq                  : STD_LOGIC_VECTOR( 31 DOWNTO 0 );     -- DMA control - assert low to enable DMA operation, high to stop DMA (for each DMA channel).
	 
	--Other signals
	SIGNAL   go                         : STD_LOGIC;
	 
	--Select signals for user's memories / reggroups
	SIGNAL   sel_reset_singlea          : STD_LOGIC;                           -- select for reset_singlea
	SIGNAL   sel_singlea_dst            : STD_LOGIC;                           -- select for singlea_dst
	 
	--FIFO SingleA
	SIGNAL   pll_mem_clk                : STD_LOGIC;
	SIGNAL   pll_write_clk              : STD_LOGIC;
	SIGNAL   pll_write_clk_pre_phy_clk  : STD_LOGIC;
	SIGNAL   pll_addr_cmd_clk           : STD_LOGIC;
	SIGNAL   pll_hr_clk                 : STD_LOGIC;
	SIGNAL   pll_p2c_read_clk           : STD_LOGIC;
	SIGNAL   pll_c2p_write_clk          : STD_LOGIC;
	SIGNAL   pll_avl_clk                : STD_LOGIC;
	SIGNAL   pll_config_clk             : STD_LOGIC;
	SIGNAL   pll_locked                 : STD_LOGIC;
	SIGNAL   afi_clk                    : STD_LOGIC;
	SIGNAL   afi_half_clk               : STD_LOGIC;
	SIGNAL   Bank_B_ready               : STD_LOGIC;                           -- 1: Memory controller is ready for use, 0: Initializing (due to reset)
	SIGNAL   data_src                   : STD_LOGIC_VECTOR( 63 DOWNTO 0 );     -- Data to the port src of FIFO singlea
	SIGNAL   singlea_flush              : STD_LOGIC;                           -- Flush FIFO data (assert high when the transfer is over)
	SIGNAL   data_dst                   : STD_LOGIC_VECTOR( 255 DOWNTO 0 );    -- Data from the port dst of FIFO singlea
	SIGNAL   wr_req_singlea             : STD_LOGIC;                           -- FIFO singlea write request signal
	SIGNAL   wr_ack_singlea             : STD_LOGIC;                           -- FIFO singlea write acknowledge signal
	SIGNAL   almost_full_singlea        : STD_LOGIC;                           -- FIFO singlea almost full signal
	SIGNAL   almost_empty_singlea       : STD_LOGIC;                           -- FIFO singlea almost empty signal
	SIGNAL   half_full_singlea          : STD_LOGIC;                           -- FIFO singlea half full signal
	SIGNAL   g_dreq_singlea             : STD_LOGIC;                           -- DMA transfer hold request from FIFO singlea
	SIGNAL   singlea_eos                : STD_LOGIC;                           -- 1: singlea port End of Stream pulse
	SIGNAL   singlea_rewind             : STD_LOGIC;                           -- 1: Start read port from the beginning of the FIFO
	 
	 
	BEGIN
		 
		 
		 
		 
		--======================================================================
		--=    The Interface entity connections (connections to the host)      =
		--======================================================================
		if_tile : tile_if
		PORT MAP  (
		 
		--Clocks & Globals
		ref_clk                      =>  ref_clk,                                  -- IN        25 MHz reference clock input pin
		clk0                         =>  clk0,                                     -- OUT       Main system clock, the max frequency is 300 MHZ
		clk                          =>  clk,                                      -- OUT       User clock, the frequency is twice/triply the frequency of clk0
		clk2                         =>  clk2,                                     -- OUT       Is an auxiliary clock that may be used as a slow emulation clock
		mem_ref_clk_int              =>  mem_ref_clk_int,                          -- OUT       Is an internal (from PLL) memory reference clock (125MHz)
		scl                          =>  scl,                                      -- INOUT     Serial clock. Used to synchronize communication to and from the I2C bus
		sda                          =>  sda,                                      -- INOUT     Serial data: Used to transfer addresses and data into and out of the I2C bus
		status_ledn( 3  DOWNTO 1 )   =>  status_ledn( 3  DOWNTO 1 ),               -- OUT       Status LEDs; 0: light on
		id( 2  DOWNTO 0 )            =>  id( 2  DOWNTO 0 ),                        -- OUT       FPGA number identification
		g_reserved( 33 DOWNTO 0 )    =>  g_reserved( 33 DOWNTO 0 ),                -- INOUT     Gidel reserved IO bus
		g_reserved_control( 99 DOWNTO 0 )  =>  g_reserved_control( 99 DOWNTO 0 ),  -- OUT       Gidel reserved control bus (out)
		 
		--PCIe connection
		pcie_refclk                  =>  pcie_refclk,                              -- IN        Reference clock for the Hard IP for PCI Express
		pcie_perst                   =>  pcie_perst,                               -- IN        Active low reset from the PCIe reset pin of the device
		pcie_rx( 7  DOWNTO 0 )       =>  pcie_rx( 7  DOWNTO 0 ),                   -- IN        Receive inputs. These signals are the serial inputs of lanes 7�0
		pcie_tx( 7  DOWNTO 0 )       =>  pcie_tx( 7  DOWNTO 0 ),                   -- OUT       Transmit outputs. These signals are the serial outputs of lanes 7�0
		 
		--Internal Bus Interface Signals
		clrn                         =>  clrn,                                     -- OUT       User Global Clear   (0: clear all)
		lclk                         =>  lclk,                                     -- OUT       Local Bus Clock
		l_wr                         =>  l_wr,                                     -- OUT       User Write Signal (1:write)
		addr_wr( 31 DOWNTO 0 )       =>  addr_wr( 31 DOWNTO 0 ),                   -- OUT       local bus address for write operations (including burst auto address increment)
		l_data_wr( 255 DOWNTO 0 )    =>  l_data_wr( 255 DOWNTO 0 ),                -- OUT       user input local data bus
		mem_ready_wr                 =>  mem_ready_wr,                             -- IN        1: end of data write transfer (memory data is valid) on rising edge of lclk
		l_rd                         =>  l_rd,                                     -- OUT       User Read Signal (0:read)
		addr_rd( 31 DOWNTO 0 )       =>  addr_rd( 31 DOWNTO 0 ),                   -- OUT       local bus address for read operations (including burst auto address increment)
		l_data_rd( 255 DOWNTO 0 )    =>  l_data_rd( 255 DOWNTO 0 ),                -- IN        data to read back from device memories
		mem_ready_rd                 =>  mem_ready_rd,                             -- IN        1: end of data read transfer (memory data is valid) on rising edge of lclk
		 
		--Interrupt Logic
		interrupt                    =>  interrupt,                                -- IN        User interrupt
		interrupt_ack                =>  interrupt_ack,                            -- OUT       User interrupt acknowledge
		 
		--DREQ Logic
		user_dreq( 31 DOWNTO 0 )     =>  user_dreq( 31 DOWNTO 0 ),                 -- IN        User DMA control for each DMA channel
		 
		--Hardware status registers (FPGA->Host)
		done                         =>  done,                                     -- IN   
		rbf_version( 7  DOWNTO 0 )   =>  rbf_version( 7  DOWNTO 0 ),               -- IN        RBF_Info[7..0]
		almost_full_dst              =>  almost_full_dst,                          -- IN        status_dst[1]
		 
		--Mode registers (Host->FPGA). Use to set hardware working modes
		go                           =>  go,                                       -- OUT  
		 
		--Select signals for user's memories / reggroups
		sel_reset_singlea            =>  sel_reset_singlea,                        -- OUT       select for reset_singlea
		sel_singlea_dst              =>  sel_singlea_dst,                          -- OUT       select for singlea_dst
		g_dreq_rd                    =>  g_dreq_singlea                            -- IN   
		);

		 
		 
		 
		--*********** START *************
		 
		--g_mp_pll_sv
		g_mp_pll_sv_cmp : g_mp_pll_sv
		PORT MAP  (
		clrn                         =>  clrn,                                     -- IN   
		mem_ref_clk                  =>  mem_ref_clk,                              -- IN   
		pll_mem_clk                  =>  pll_mem_clk,                              -- OUT  
		pll_write_clk                =>  pll_write_clk,                            -- OUT  
		pll_write_clk_pre_phy_clk    =>  pll_write_clk_pre_phy_clk,                -- OUT  
		pll_addr_cmd_clk             =>  pll_addr_cmd_clk,                         -- OUT  
		pll_hr_clk                   =>  pll_hr_clk,                               -- OUT  
		pll_p2c_read_clk             =>  pll_p2c_read_clk,                         -- OUT  
		pll_c2p_write_clk            =>  pll_c2p_write_clk,                        -- OUT  
		pll_avl_clk                  =>  pll_avl_clk,                              -- OUT  
		pll_config_clk               =>  pll_config_clk,                           -- OUT  
		pll_locked                   =>  pll_locked,                               -- OUT  
		afi_clk                      =>  afi_clk,                                  -- OUT  
		afi_half_clk                 =>  afi_half_clk                              -- OUT  
		);

		 
		 
		 
		 
		--======================================================================
		--=                   User's entities' connections                     =
		--======================================================================
		 
		 
		--user
		 
		user_cmp : user
		PORT MAP  (
		clrn                         =>  clrn,                                     -- IN   
		clk0                         =>  clk0,                                     -- IN   
		go                           =>  go,                                       -- IN   
		done                         =>  done,                                     -- OUT  
		Bank_B_ready                 =>  Bank_B_ready,                             -- IN        1: Memory controller is ready for use, 0: Initializing (due to reset)
		data_src                     =>  data_src,                                 -- OUT       Data to the port src of FIFO singlea
		wr_req_singlea               =>  wr_req_singlea,                           -- OUT       FIFO singlea write request signal
		wr_ack_singlea               =>  wr_ack_singlea,                           -- IN        FIFO singlea write acknowledge signal
		singlea_eos                  =>  singlea_eos,                              -- IN        1: singlea port End of Stream pulse
		singlea_flush                =>  singlea_flush,                            -- OUT       Flush FIFO data (assert high when the transfer is over)
		singlea_rewind               =>  singlea_rewind                            -- OUT       1: Start read port from the beginning of the FIFO
		);

		 
		 
		 
		--*********** FINISH *************
		 
		 
		--======================================================================
		--=                   SDRAM controllers' connections                   =
		--======================================================================
		 
		--======================================================================
		--=                         IC_1_Bank_B_Ctrl                           =
		--======================================================================
		 
		 
		IC_1_Bank_B_Ctrl_cmp : IC_1_Bank_B_Ctrl
		PORT MAP  (
		 
		--Global MultiPort Connections
		clrn                         =>  clrn,                                     -- IN   
		ref_clk                      =>  mem_ref_clk,                              -- IN   
		pll_mem_clk                  =>  pll_mem_clk,                              -- IN   
		pll_write_clk                =>  pll_write_clk,                            -- IN   
		pll_write_clk_pre_phy_clk    =>  pll_write_clk_pre_phy_clk,                -- IN   
		pll_addr_cmd_clk             =>  pll_addr_cmd_clk,                         -- IN   
		pll_hr_clk                   =>  pll_hr_clk,                               -- IN   
		pll_p2c_read_clk             =>  pll_p2c_read_clk,                         -- IN   
		pll_c2p_write_clk            =>  pll_c2p_write_clk,                        -- IN   
		pll_avl_clk                  =>  pll_avl_clk,                              -- IN   
		pll_config_clk               =>  pll_config_clk,                           -- IN   
		pll_locked                   =>  pll_locked,                               -- IN   
		afi_clk                      =>  afi_clk,                                  -- IN   
		afi_half_clk                 =>  afi_half_clk,                             -- IN   
		g_reserved_control( 99 DOWNTO 0 )  =>  g_reserved_control( 99 DOWNTO 0 ),  -- IN   
		ready                        =>  Bank_B_ready,                             -- OUT  
		 
		--SDRAM Connections
		data( 63 DOWNTO 0 )          =>  dq_b( 63 DOWNTO 0 ),                      -- OUT  
		addr( 15 DOWNTO 0 )          =>  addr_b( 15 DOWNTO 0 ),                    -- OUT  
		dqm( 7  DOWNTO 0 )           =>  dqm_b( 7  DOWNTO 0 ),                     -- OUT  
		dqs( 7  DOWNTO 0 )           =>  dqs_b( 7  DOWNTO 0 ),                     -- OUT  
		dqsn( 7  DOWNTO 0 )          =>  dqsn_b( 7  DOWNTO 0 ),                    -- OUT  
		ba( 2  DOWNTO 0 )            =>  ba_b( 2  DOWNTO 0 ),                      -- OUT  
		cs_bus( 1  DOWNTO 0 )        =>  cs_b( 1  DOWNTO 0 ),                      -- OUT  
		ce( 1  DOWNTO 0 )            =>  cke_b( 1  DOWNTO 0 ),                     -- OUT  
		ras                          =>  ras_b,                                    -- OUT  
		cas                          =>  cas_b,                                    -- OUT  
		we                           =>  we_b,                                     -- OUT  
		odt( 1  DOWNTO 0 )           =>  odt_b( 1  DOWNTO 0 ),                     -- OUT  
		ck( 1  DOWNTO 0 )            =>  ck_b( 1  DOWNTO 0 ),                      -- OUT  
		ckn( 1  DOWNTO 0 )           =>  ckn_b( 1  DOWNTO 0 ),                     -- OUT  
		oct_rzqin                    =>  rzq_b,                                    -- OUT  
		event_in                     =>  event_b,                                  -- OUT  
		mem_reset_n                  =>  resetn_b,                                 -- OUT  
		 
		--Port src of FIFO singlea Connections
		clk_src                      =>  clk0,                                     -- IN   
		data_src( 63 DOWNTO 0 )      =>  data_src( 63 DOWNTO 0 ),                  -- IN   
		singlea_flush                =>  singlea_flush,                            -- IN   
		 
		--Port dst of FIFO singlea Connections
		clk_dst                      =>  lclk,                                     -- IN   
		data_dst( 255 DOWNTO 0 )     =>  data_dst( 255 DOWNTO 0 ),                 -- OUT  
		singlea_almost_full_dst      =>  almost_full_dst,                          -- OUT  
		 
		--FIFO singlea Connections
		reset_singlea                =>  sel_reset_singlea,                        -- IN   
		lclk                         =>  lclk,                                     -- IN   
		sel_singlea                  =>  sel_singlea_dst,                          -- IN   
		wr_req_singlea               =>  wr_req_singlea,                           -- IN   
		wr_ack_singlea               =>  wr_ack_singlea,                           -- OUT  
		almost_full_singlea          =>  almost_full_singlea,                      -- OUT  
		almost_empty_singlea         =>  almost_empty_singlea,                     -- OUT  
		half_full_singlea            =>  half_full_singlea,                        -- OUT  
		g_dreq_singlea               =>  g_dreq_singlea,                           -- OUT  
		singlea_eos                  =>  singlea_eos,                              -- OUT  
		singlea_rewind               =>  singlea_rewind                            -- IN   
		);

		 
		 
		rbf_version(7 DOWNTO 0)    <=    RBF_VERSION_VAL;  
		 
		 
		--======================================================================
		--=                Default Values of Board Connections                 =
		--======================================================================
		 
		--DDR Block C Connections
		addr_c                       <=  ( others => '0' );
		ba_c                         <=  ( others => '0' );
		cas_c                        <=  '1';
		cke_c                        <=  ( others => '0' );
		ck_c                         <=  ( others => 'Z' );
		ckn_c                        <=  ( others => 'Z' );
		cs_c                         <=  ( others => '1' );
		dq_c                         <=  ( others => 'Z' );
		dqm_c                        <=  ( others => '0' );
		dqs_c                        <=  ( others => 'Z' );
		dqsn_c                       <=  ( others => 'Z' );
		we_c                         <=  '0';
		ras_c                        <=  '1';
		odt_c                        <=  ( others => '0' );
		resetn_c                     <=  '0';
		 
		--DDR Block D Connections
		dq_d                         <=  ( others => 'Z' );
		ldn_d                        <=  '1';
		bwsn_d                       <=  ( others => '0' );
		r_wn_d                       <=  '0';
		k_d                          <=  '0';
		addr_d                       <=  ( others => '0' );
		 
		--DDR Block D Connections
		dq_e                         <=  ( others => 'Z' );
		ldn_e                        <=  '1';
		bwsn_e                       <=  ( others => '0' );
		r_wn_e                       <=  '0';
		k_e                          <=  '0';
		addr_e                       <=  ( others => '0' );
		 
		--User's buses
		 
		mem_ready_wr                 <=  '1';                                      -- '1'   NO WAIT STATES, put '0' when you want to add wait states
		 
		mem_ready_rd                 <=  '1';                                      -- '1'   NO WAIT STATES, put '0' when you want to add wait states
		l_data_rd( 31 DOWNTO 0 )     <= data_dst( 31 DOWNTO 0 )   WHEN   sel_singlea_dst  =  '1'   ELSE
		                              ( others => '0' );
		 
		l_data_rd( 255 DOWNTO 32 )   <= data_dst( 255 DOWNTO 32 )   WHEN   sel_singlea_dst  =  '1'   ELSE
		                              ( others => '0' );
		 
		interrupt                    <=  '1';                                      -- Interrupt control - assert low to send interrupt to SoftWare, when interrupt_ack is high.
		user_dreq                    <=  ( others => '0' );                        -- DMA control - assert low to enable DMA operation, high to stop DMA (for each DMA channel).
		ledn                         <=  ( others => 'Z' );
		 
		--1G PHY I/O's (Connections to on board PHY)
		phy_mdio                     <=  'Z';
		phy_mdc                      <=  '0';
		phy_resetn                   <=  '0';
		phy_tx_ctrl                  <=  '0';
		phy_tx_clk                   <=  '0';
		phy_txd                      <=  ( others => '0' );
		 
		--SFP A
		sfp_link_ledn_a              <=  'Z';
		sfp_trafic_ledn_a            <=  'Z';
		 
		--SFP B
		sfp_link_ledn_b              <=  'Z';
		sfp_trafic_ledn_b            <=  'Z';
		 
		--L(J4) connector I/O's
		l                            <=  ( others => 'Z' );
		l_io                         <=  ( others => 'Z' );
		clk_out                      <=  ( others => '0' );
		 
		--External(J3) connector I/O's
		j3_ext_io                    <=  ( others => 'Z' );
		j3_ext_io_dir                <=  ( others => '0' );                        -- Bit-0 sets direction for ext_io[7:0] and bit-1 for ext_io[11:8]. (ext_io_dir=0: Inputs, ext_io_dir=1: Outputs)
		 
		 
	END  tile_arch;
